class base;
randc bit in0;
randc bit in1;
randc bit sel;
bit out;
endclass
