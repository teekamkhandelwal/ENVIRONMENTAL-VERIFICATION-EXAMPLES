
`ifndef __dff_base__
`define __dff_base__

class d_pkt;
 rand bit d;
      bit q;
      bit rst;
endclass

`endif
