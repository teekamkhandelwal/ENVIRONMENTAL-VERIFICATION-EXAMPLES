`ifndef __dff_cfg__
`define __dff_cfg__

class d_cfg;
  int num_txn;
end

`endif
